module router_sync(input clock,resetn,detect_add,write_enb_reg,full_0,full_1,full_2,empty_0,empty_1,empty_2,read_enb_0,read_enb_1,read_enb_2,
                                   input [1:0] data_in,
                                   output reg [2:0] write_enb,
                                   output reg fifo_full,soft_reset_0,soft_reset_1,soft_reset_2,
                                   output vld_out_0,vld_out_1,vld_out_2);

reg [1:0] temp;
reg [4:0] count0,count1,count2;

always@(posedge clock)
        begin
                if(~resetn)
                        begin
                                temp <= 2'b10;
                        end
                else if(detect_add)
                        temp <= data_in;
        end

always@(*)
        begin
                if(write_enb_reg)
                        begin
                                case(temp)
                                        2'b00: write_enb <= 3'b001;
                                        2'b01: write_enb <= 3'b010;
                                        2'b10: write_enb <= 3'b100;
                                  default: write_enb <= 3'b000;
                                endcase
                        end
                else
                        write_enb <= 3'b000;
        end
always@(posedge clock or full_0 or full_1 or full_2)                            //because for pkt 14 when full_2 is high fifo_full is high on next posedge
        begin
                if((full_0 == 1'b1) || (full_1 == 1'b1) || (full_2 == 1'b1))
                        begin
                                case(temp)
                                        2'b00: fifo_full <= full_0;
                                        2'b01: fifo_full <= full_1;
                                        2'b10: fifo_full <= full_2;
                                        default: fifo_full <= full_0;
                                endcase
                        end
                else
                        fifo_full <= 1'd0;

        end


always@(posedge clock)
        begin
                if(~resetn)
                        begin
                                count0 <= 5'd0;
                                soft_reset_0 <= 1'b0;
                        end
                else
                begin
                        if(vld_out_0)
                                begin
                                        if(~read_enb_0)
                                                begin
                                                        if(count0 == 5'd30)
                                                                begin
                                                                        soft_reset_0 <= 1'b1;
                                                                        count0 <= 5'd0;
                                                                end
 else
                                                                begin
                                                                        count0 <= count0 + 5'd1;
                                                                        soft_reset_0 <= 1'b0;
                                                                end
                                                end
                                        else
                                        count0 <= 5'd0;
                                end
                end
        end


always@(posedge clock)
        begin
                if(~resetn)
                        begin
                                count1 <= 5'd0;
                                soft_reset_1 <= 1'b0;
                        end
                else
                begin
                        if(vld_out_1)
                                begin
                                        if(~read_enb_1)
                                                begin
                                                        if(count1 == 5'd30)
                                                                begin
                                                                        soft_reset_1 <= 1'b1;
                                                                        count1 <= 5'd0;
                                                                end
                                                        else
                                                                begin
                                                                        count1 <= count1 + 5'd1;
                                                                        soft_reset_1 <= 1'b0;
                                                                end
                                                end
  else
                                        count1 <= 5'd0;
                                end

                end
        end

always@(posedge clock)
        begin
                if(~resetn)
                        begin
                                count2 <= 5'd0;
                                soft_reset_2 <= 1'b0;
                        end
                else
                begin
                        if(vld_out_2)
                                begin
                                        if(~read_enb_2)
                                                begin
                                                        if(count2 == 5'd30)
                                                                begin
                                                                        soft_reset_2 <= 1'b1;
                                                                        count2 <= 5'd0;
                                                                end
                                                        else
                                                                begin
                                                                        count2 <= count2 + 5'd1;
                                                                        soft_reset_2 <= 1'b0;
                                                                end
                                                end
                                        else
                                        count2 <= 5'd0;
                                end

                end
        end


assign vld_out_0 = ~empty_0;
assign vld_out_1 = ~empty_1;
assign vld_out_2 = ~empty_2;

endmodule